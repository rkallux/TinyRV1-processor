//========================================================================
// ImmGen_RTL-test
//========================================================================

`include "ece2300-test.v"
`include "ImmGen_RTL.v"

module Top();

  //----------------------------------------------------------------------
  // Setup
  //----------------------------------------------------------------------

  // verilator lint_off UNUSED
  logic clk;
  logic reset;
  // verilator lint_on UNUSED

  ece2300_TestUtils t( .* );

  //----------------------------------------------------------------------
  // Instantiate design under test
  //----------------------------------------------------------------------

  logic [31:0] dut_inst;
  logic  [1:0] dut_imm_type;
  logic [31:0] dut_imm;

  ImmGen_RTL dut
  (
    .inst     (dut_inst),
    .imm_type (dut_imm_type),
    .imm      (dut_imm)
  );

  //----------------------------------------------------------------------
  // check
  //----------------------------------------------------------------------
  // All tasks start at #1 after the rising edge of the clock. So we
  // write the inputs #1 after the rising edge, and check the outputs #1
  // before the next rising edge.

  task check
  (
    input logic [31:0] inst,
    input logic  [1:0] imm_type,
    input logic [31:0] imm
  );
    if ( !t.failed ) begin

      dut_inst     = inst;
      dut_imm_type = imm_type;

      #8;

      if ( t.n != 0 ) begin
        $display( "%3d: %h %d > %h", t.cycles,
                  dut_inst, dut_imm_type, dut_imm );
      end

      `ECE2300_CHECK_EQ( dut_imm, imm );

      #2;

    end
  endtask

  //----------------------------------------------------------------------
  // test_case_1_basic
  //----------------------------------------------------------------------

  task test_case_1_basic();
    t.test_case_begin( "test_case_1_basic" );

    //     inst           imm_type imm
    check( 32'h0000_0000, 0,       32'h0000_0000 );
    check( 32'h0000_0000, 1,       32'h0000_0000 );
    check( 32'h0000_0000, 2,       32'h0000_0000 );
    check( 32'h0000_0000, 3,       32'h0000_0000 );

  endtask

  //----------------------------------------------------------------------
  // test_case_2_directed_i_type
  //----------------------------------------------------------------------

  task test_case_2_directed_i_type();
    t.test_case_begin( "test_case_2_directed_i_type" );

    //         **** **** ****                                                           **** **** ****
    check( 32'b0000_0000_0000_0000_0000_0000_0000_0000, 0, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0000_0001_0000_0000_0000_0000_0000, 0, 32'b0000_0000_0000_0000_0000_0000_0000_0001 );
    check( 32'b0101_0101_0101_0000_0000_0000_0000_0000, 0, 32'b0000_0000_0000_0000_0000_0101_0101_0101 );
    check( 32'b0110_1001_1111_0000_0000_0000_0000_0000, 0, 32'b0000_0000_0000_0000_0000_0110_1001_1111 );
    check( 32'b1000_0000_0000_0000_0000_0000_0000_0000, 0, 32'b1111_1111_1111_1111_1111_1000_0000_0000 );

    check( 32'b0000_0000_0000_1111_1111_1111_1111_1111, 0, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0000_0001_1111_1111_1111_1111_1111, 0, 32'b0000_0000_0000_0000_0000_0000_0000_0001 );
    check( 32'b0101_0101_0101_1111_1111_1111_1111_1111, 0, 32'b0000_0000_0000_0000_0000_0101_0101_0101 );
    check( 32'b0110_1001_1111_1111_1111_1111_1111_1111, 0, 32'b0000_0000_0000_0000_0000_0110_1001_1111 );
    check( 32'b1000_0000_0000_1111_1111_1111_1111_1111, 0, 32'b1111_1111_1111_1111_1111_1000_0000_0000 );

  endtask

  //----------------------------------------------------------------------
  // test_case_3_directed_s_type
  //----------------------------------------------------------------------

  task test_case_3_directed_s_type();
    t.test_case_begin( "test_case_3_directed_s_type" );

    //         **** ***                 **** *                                          **** **** ****
    check( 32'b0000_0000_0000_0000_0000_0000_0000_0000, 1, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0000_0000_0000_0000_0000_1000_0000, 1, 32'b0000_0000_0000_0000_0000_0000_0000_0001 );
    check( 32'b0010_1010_0000_0000_0000_1010_1000_0000, 1, 32'b0000_0000_0000_0000_0000_0010_1011_0101 );
    check( 32'b0110_1010_0000_0000_0000_1111_1000_0000, 1, 32'b0000_0000_0000_0000_0000_0110_1011_1111 );
    check( 32'b1000_0000_0000_0000_0000_0000_0000_0000, 1, 32'b1111_1111_1111_1111_1111_1000_0000_0000 );

    check( 32'b0000_0001_1111_1111_1111_0000_0111_1111, 1, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0001_1111_1111_1111_0000_1111_1111, 1, 32'b0000_0000_0000_0000_0000_0000_0000_0001 );
    check( 32'b0010_1011_1111_1111_1111_1010_1111_1111, 1, 32'b0000_0000_0000_0000_0000_0010_1011_0101 );
    check( 32'b0110_1011_1111_1111_1111_1111_1111_1111, 1, 32'b0000_0000_0000_0000_0000_0110_1011_1111 );
    check( 32'b1000_0001_1111_1111_1111_0000_0111_1111, 1, 32'b1111_1111_1111_1111_1111_1000_0000_0000 );

  endtask

  //----------------------------------------------------------------------
  // test_case_4_directed_j_type
  //----------------------------------------------------------------------

  task test_case_4_directed_j_type();
    t.test_case_begin( "test_case_4_directed_j_type" );

    //         abbb bbbb bbbc dddd dddd                                     a dddd dddd cbbb bbbb bbb0
    check( 32'b0000_0000_0000_0000_0000_0000_0000_0000, 2, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0000_0010_0000_0000_0000_0000_0000, 2, 32'b0000_0000_0000_0000_0000_0000_0000_0010 );
    check( 32'b0010_1010_1011_1010_1010_0000_0000_0000, 2, 32'b0000_0000_0000_1010_1010_1010_1010_1010 );
    check( 32'b1000_0000_0000_0000_0000_0000_0000_0000, 2, 32'b1111_1111_1111_0000_0000_0000_0000_0000 );

    check( 32'b0000_0000_0000_0000_0000_1111_1111_1111, 2, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0000_0010_0000_0000_1111_1111_1111, 2, 32'b0000_0000_0000_0000_0000_0000_0000_0010 );
    check( 32'b0010_1010_1011_1010_1010_1111_1111_1111, 2, 32'b0000_0000_0000_1010_1010_1010_1010_1010 );
    check( 32'b1000_0000_0000_0000_0000_1111_1111_1111, 2, 32'b1111_1111_1111_0000_0000_0000_0000_0000 );

  endtask

  //----------------------------------------------------------------------
  // test_case_5_directed_b_type
  //----------------------------------------------------------------------

  task test_case_5_directed_b_type();
    t.test_case_begin( "test_case_5_directed_b_type" );

    //         abbb bbb                 dddd c                                        a cbbb bbbd ddd0
    check( 32'b0000_0000_0000_0000_0000_0000_0000_0000, 3, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0000_0000_0000_0000_0001_0000_0000, 3, 32'b0000_0000_0000_0000_0000_0000_0000_0010 );
    check( 32'b0010_1010_0000_0000_0000_0101_1000_0000, 3, 32'b0000_0000_0000_0000_0000_1010_1010_1010 );
    check( 32'b1000_0000_0000_0000_0000_0000_0000_0000, 3, 32'b1111_1111_1111_1111_1111_0000_0000_0000 );

    check( 32'b0000_0001_1111_1111_1111_0000_0111_1111, 3, 32'b0000_0000_0000_0000_0000_0000_0000_0000 );
    check( 32'b0000_0001_1111_1111_1111_0001_0111_1111, 3, 32'b0000_0000_0000_0000_0000_0000_0000_0010 );
    check( 32'b0010_1011_1111_1111_1111_0101_1111_1111, 3, 32'b0000_0000_0000_0000_0000_1010_1010_1010 );
    check( 32'b1000_0001_1111_1111_1111_0000_0111_1111, 3, 32'b1111_1111_1111_1111_1111_0000_0000_0000 );

  endtask

  //----------------------------------------------------------------------
  // main
  //----------------------------------------------------------------------

  initial begin
    t.test_bench_begin( `__FILE__ );

    if ((t.n <= 0) || (t.n == 1)) test_case_1_basic();
    if ((t.n <= 0) || (t.n == 2)) test_case_2_directed_i_type();
    if ((t.n <= 0) || (t.n == 3)) test_case_3_directed_s_type();
    if ((t.n <= 0) || (t.n == 4)) test_case_4_directed_j_type();
    if ((t.n <= 0) || (t.n == 5)) test_case_5_directed_b_type();

    t.test_bench_end();
  end

endmodule

